    `include "uart_trans.sv"
    `include "uart_agent_cfg.sv"
    
    `include "uart_sequence.sv"
    `include "uart_sequencer.sv"
    
    `include "uart_mon.sv"
    `include "uart_driver.sv"

    `include "uart_agent.sv"
