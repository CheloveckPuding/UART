`timescale 1ns/10ps
interface uart_intf;
  
  logic rx;
  logic tx;


endinterface
