    `include "uart_trans.svh"
    
    `include "uart_sequence.svh"
    
    `include "uart_mon.svh"
    `include "uart_driver.svh"

    `include "uart_agent.svh"
